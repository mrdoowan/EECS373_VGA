`timescale 1ns / 1ps 
////////////////////////////////////////////////////////////////////////////////// 
//  
// Source Code is inspired from: 
// https://www.element14.com/community/thread/23394/l/draw-vga-color-bars-with-fpga-in-verilog?displayFullThread=true 
// Code has been modified to meet the needs for the EECS 373 Final Project at Winter 2016
// Coded by: Steven Duan 
// 
////////////////////////////////////////////////////////////////////////////////// 

// ------------------------------------------------------ 
// MAIN MODULE 
// ------------------------------------------------------ 

module eecs373_VGA( 
	 input wire clk,           //master clock = 50MHz 
	 input wire clr, 	         //Reset SW17, for Clock Divider and VGA
	 input wire KEY3,         	//Increment Player 1 points 
	 input wire KEY2,         	//Increment Player 2 points
	 input wire KEY1,				//Change colors
	 input wire KEY0,				//Resets Player score 
	 input wire SCLK,				//Clock from SPI device
	 input wire MOSI,				//Master out, Slave in data
	 input wire SSEL,				//Slave select
	 input wire SW0,				//To switch between KEY increment / SPI 
	 input wire SW1,				//To switch between P1 and P2 for colors
	 output reg [15:0] byte_data_received, // SPI data from Master
	 output wire GPIO1,
	 output wire VGA_CLK,     	//VGA display clock interconnect (25MHz) 
	 output wire n_sync,       //Determines if sync-on-green is used. Set to '0' 
	 output wire n_blank,      //Determines if direct blanking is used. Set to '1' 
	 output wire [7:0] red,    //red vga output - 8 bits 
	 output wire [7:0] green,  //green vga output - 8 bits 
	 output wire [7:0] blue,   //blue vga output - 8 bits 
	 output wire hsync,        //horizontal sync out 
	 output wire vsync,        //vertical sync out 
	 output wire [6:0] HEX7,  	//P1 score on 7seg 
	 output wire [6:0] HEX6,  	//P1 score on 7seg 
	 output wire [6:0] HEX5,  	//P2 score on 7seg 
	 output wire [6:0] HEX4   	//P2 score on 7seg 
	 ); 
	  
	  // Assigning respective values for VGA
	 assign n_sync = 0; 
	 assign n_blank = 1; 
		
	 // Only purpose is to see the clock.
	 assign GPIO1 = VGA_CLK;
	 
	 // Debounced Switches 
	 wire reset_deb; 
	 wire KEY2_deb; 
	 wire KEY3_deb; 
	 wire KEY1_deb;
	  
		debouncer d0( 
		  .clk(clk), 
		  .PB(KEY0), 
		  .PB_state(reset_deb) 
		); 
		// Detect reset falling edge
		reg [2:0] reset_r;
		always @(posedge clk) reset_r <= {reset_r[1:0], reset_deb};
		wire Reset_fallingedge = (reset_r[2:1] == 2'b10);
		
		debouncer d3( 
		  .clk(clk), 
		  .PB(KEY3), 
		  .PB_state(KEY3_deb) 
		); 
		// Detect KEY3 falling edge
		reg [2:0] KEY3_r;
		always @(posedge clk) KEY3_r <= {KEY3_r[1:0], KEY3_deb};
		wire KEY3_fallingedge = (KEY3_r[2:1] == 2'b10);
		
		debouncer d2( 
		  .clk(clk), 
		  .PB(KEY2), 
		  .PB_state(KEY2_deb) 
		); 
		// Detect KEY2 falling edge
		reg [2:0] KEY2_r;
		always @(posedge clk) KEY2_r <= {KEY2_r[1:0], KEY2_deb};
		wire KEY2_fallingedge = (KEY2_r[2:1] == 2'b10);
	
		
		debouncer d1( 
		  .clk(clk), 
		  .PB(KEY1), 
		  .PB_state(KEY1_deb) 
		); 
		// Detect KEY1 falling edge
		reg [2:0] KEY1_r;
		always @(posedge clk) KEY1_r <= {KEY1_r[1:0], KEY1_deb};
		wire KEY1_fallingedge = (KEY1_r[2:1] == 2'b10);
		
		// Generate pixel clock by using a clock divider 
		clockdiv U1( 
		  .clk(clk), 
		  .reset(clr), 
		  .VGA_CLK(VGA_CLK) 
		  ); 
		
	  //----------------------------------------------------
	  // (BELOW) SPI Module
	  // (Credit goes to http://www.fpga4fun.com/SPI2.html)
	  //----------------------------------------------------
	  
		// sync SCLK to the FPGA Clock
		reg [2:0] SCLKr;
		always @(posedge clk) SCLKr <= {SCLKr[1:0], SCLK};
		wire SCLK_risingedge = (SCLKr[2:1] == 2'b01); // Detect SPI clk rising edge
		wire SCLK_fallingedge = (SCLKr[2:1] == 2'b10); // Detect SPI clk falling edge
		
		// sync SSEL to the FPGA Clock
		reg [2:0] SSELr;
		always @(posedge clk) SSELr <= {SSELr[1:0], SSEL};
		wire SSEL_active = ~SSELr[1];			// SSEL is active low
		// Do not need to use SSEL_message since we are not transmitting
		
		// sync MOSI to the FPGA Clock
		reg [1:0] MOSIr;
		always @(posedge clk) MOSIr <= {MOSIr[0], MOSI};
		wire MOSI_data = MOSIr[1];
		
		// SPI messages being sent is being done in a 16-bit format
		reg [3:0] bitcount;	// Counts up to 16
		reg data_received; 	// T/F if data was received
		
		always @(posedge clk)
		begin
			if (~SSEL_active)
				bitcount <= 0;
			else if (SCLK_risingedge)
			begin
				bitcount <= bitcount + 1;
				// Left shift register on the byte_data received
				byte_data_received <= {byte_data_received[14:0], MOSI_data};
			end
		end
		
		// Just to check if the full 2 bytes was received
		always @(posedge clk) data_received = SSEL_active && SCLK_risingedge && (bitcount == 15);
		
	  //----------------------------------------------------
	  // (ABOVE) SPI Module
	  //----------------------------------------------------
	  
	  // 1st Byte
	  // This represents that Player 1/2 score needs to be updated!
	  // byte_data_received[15] = Player 1 (0) / Player 2 (1)
	  // byte_data_received[14:8] = Points
	  // 2nd Byte
	  // byte_data_received[7:0] = State of RGB
	  
	  //-----------------------------------------------------
	  // (BELOW) Color Switching
	  //-----------------------------------------------------
	  
	  parameter BLUE1 = 3'b000;
	  parameter RED1 = 3'b001;
	  parameter RED2 = 3'b000;
	  parameter BLUE2 = 3'b001;
	  parameter GREEN = 3'b010;
	  parameter YELLOW = 3'b011;
	  parameter PURPLE = 3'b100;
	  parameter CYAN = 3'b101;
	  
	  reg [7:0] state1;
	  reg [7:0] state2;
	  
	  // Cycle around the states
	  always @(posedge clk)
	  begin
			if (~byte_data_received[15] && data_received)
				state1 <= byte_data_received[7:0];
			else if (byte_data_received[15] && data_received)
				state2 <= byte_data_received[7:0];
	  end
	  
	  // To hold colors: [23:16] <= Red, [15:8] <= Green, [7:0] Blue
	  reg [23:0] color1;
	  reg [23:0] color2;
	  
	  // Combinational output
	  always @*
	  begin
			case(state1)	  //24'bRRRRRRRRGGGGGGGGBBBBBBBB
			RED1:		color1 <= 24'b111111110000000000000000;
			GREEN:	color1 <= 24'b000000001100110000000000;
			YELLOW:	color1 <= 24'b111111111111111100000000;
			PURPLE:	color1 <= 24'b110011000000000011001100;
			CYAN:		color1 <= 24'b000000001111111111111111;
			default:	color1 <= 24'b000000001000000011111111;
			endcase
	  end
	  
	  always @*
	  begin
			case(state2)	  //24'bRRRRRRRRGGGGGGGGBBBBBBBB
			BLUE2:	color2 <= 24'b000000001000000011111111;
			GREEN:	color2 <= 24'b000000001100110000000000;
			YELLOW:	color2 <= 24'b111111111111111100000000;
			PURPLE:	color2 <= 24'b110011000000000011001100;
			CYAN:		color2 <= 24'b000000001111111111111111;
			default:	color2 <= 24'b111111110000000000000000;
			endcase
	  end
	  
	  //-----------------------------------------------------
	  // (ABOVE) Color Switching
	  //-----------------------------------------------------

	  //-----------------------------------------------------
	  // (BELOW) Logic for Incrementing Points
	  //-----------------------------------------------------
	  
	  // Counter for how many points
	  reg [6:0] P1_points; 
	  reg [6:0] P2_points;
	  
	  // There are two different modes on how the Points are being handled
	  // ~SW0 (when the switch is low) is when points are from the SPI
	  // SW0 (when the switch is high) is when points are incremented by Key Button
	  always @(posedge clk)
	  begin
		  // Data from SPI
		  if (~byte_data_received[15] && ~SW0 && data_received)
		  begin
			  P1_points <= byte_data_received[14:8];
		  end
		  else if (byte_data_received[15] && ~SW0 && data_received)
		  begin
			  P2_points <= byte_data_received[14:8];
		  end
		  // Data from Key Button
		  else if (KEY3_fallingedge && SW0)
		  begin
			  if (P1_points >= 99) P1_points <= 99; 
			  else P1_points <= P1_points + 1; 
		  end
		  else if (KEY2_fallingedge && SW0)
		  begin
			  if (P2_points >= 99) P2_points <= 99; 
			  else P2_points <= P2_points + 1; 
		  end
		  // Resets the points back to zero
		  else if (Reset_fallingedge)
		  begin
			  P1_points <= 0;
			  P2_points <= 0;
		  end
	  end
		
	  //-----------------------------------------------------
	  // (ABOVE) Logic for Incrementing Points
	  //-----------------------------------------------------	
	
	  // Combinational Logic for Output 
	  wire [3:0] single1 = P1_points % 10; 
	  wire [3:0] single2 = P2_points % 10;
	
	  // Display points on 7 Segment Hex. 
	  display_hex seg7( 
			 .P1(P1_points), 
			 .P2(P2_points), 
			 .S1(single1), 
			 .S2(single2), 
			 .HEX7(HEX7), 
			 .HEX6(HEX6), 
			 .HEX5(HEX5), 
			 .HEX4(HEX4) 
			 ); 
		
	  // ---------------------------------------- 
	  // VGA Display 
	  // ---------------------------------------- 
	 vga640x480 U3( 
			.VGA_CLK(VGA_CLK), 
			.P1(P1_points), 
			.P2(P2_points), 
			.S1(single1), 
			.S2(single2),
			.color1(color1),
			.color2(color2),
			.reset(clr), 
			.hsync(hsync), 
			.vsync(vsync), 
			.red(red), 
			.green(green), 
			.blue(blue) 
			); 
	  
endmodule 

// ------------------------------------------------------ 
// ------------------------------------------------------ 
// ------------------------------------------------------ 
// ADDITIONAL MODULES. MAIN MODULE ABOVE 
// ------------------------------------------------------ 
// ------------------------------------------------------ 
// ------------------------------------------------------ 

// ------------------------------------------------------ 
// Submodule: Clock Divider 
// ------------------------------------------------------ 

module clockdiv( 
	 input wire clk,        //master clock: 50MHz 
	 input wire reset,      //SW17 button reset 
	 output wire VGA_CLK       //pixel clock: 25MHz 
	 ); 

	 // 17-bit counter variable 
	 reg [31:0] counter; 

	 // Clock divider -- 
	 // Used to divide the clock from 50MHz 
	 always @(posedge clk) 
	 begin 
		// reset condition 
		  if (reset) 
				counter <= 0; 
		  else 
				counter <= counter + 1; 
	 end 
		
	 // 50Mhz ÷ 2^1 = 25MHz 
	 assign VGA_CLK = counter[0]; 

endmodule 

// ------------------------------------------------------ 
// Submodule: Hex Display 
// ------------------------------------------------------ 

module display_hex( 
	 input wire [6:0] P1, 
	 input wire [6:0] P2, 
	 input wire [3:0] S1, 
	 input wire [3:0] S2, 
	 output reg [6:0] HEX7, 
	 output reg [6:0] HEX6, 
	 output reg [6:0] HEX5, 
	 output reg [6:0] HEX4 
	 ); 

	 parameter n0 = 7'b1000000; 
	 parameter n1 = 7'b1111001; 
	 parameter n2 = 7'b0100100; 
	 parameter n3 = 7'b0110000; 
	 parameter n4 = 7'b0011001; 
	 parameter n5 = 7'b0010010; 
	 parameter n6 = 7'b0000010; 
	 parameter n7 = 7'b1111000; 
	 parameter n8 = 7'b0000000; 
	 parameter n9 = 7'b0011000; 
	  
	 always @* 
	 begin 
		  // Player 1 display on HEX7, HEX6 
		  // HEX7 
		  begin 
				if (P1 >= 0 && P1 < 10) HEX7 <= n0;  
				else if (P1 >= 10 && P1 < 20) HEX7 <= n1; 
				else if (P1 >= 20 && P1 < 30) HEX7 <= n2; 
				else if (P1 >= 30 && P1 < 40) HEX7 <= n3; 
				else if (P1 >= 40 && P1 < 50) HEX7 <= n4; 
				else if (P1 >= 50 && P1 < 60) HEX7 <= n5; 
				else if (P1 >= 60 && P1 < 70) HEX7 <= n6; 
				else if (P1 >= 70 && P1 < 80) HEX7 <= n7; 
				else if (P1 >= 80 && P1 < 90) HEX7 <= n8; 
				else HEX7 <= n9; 
		  end 
		  // HEX6 
		  begin 
				if (S1 == 0) HEX6 <= n0; 
				else if (S1 == 1) HEX6 <= n1; 
				else if (S1 == 2) HEX6 <= n2; 
				else if (S1 == 3) HEX6 <= n3; 
				else if (S1 == 4) HEX6 <= n4; 
				else if (S1 == 5) HEX6 <= n5; 
				else if (S1 == 6) HEX6 <= n6; 
				else if (S1 == 7) HEX6 <= n7; 
				else if (S1 == 8) HEX6 <= n8; 
				else HEX6 <= n9; 
		  end 
		  // Player 2 display on HEX5, HEX4 
		  // HEX5 
		  begin 
				if (P2 >= 0 && P2 < 10) HEX5 <= n0;  
				else if (P2 >= 10 && P2 < 20) HEX5 <= n1; 
				else if (P2 >= 20 && P2 < 30) HEX5 <= n2; 
				else if (P2 >= 30 && P2 < 40) HEX5 <= n3; 
				else if (P2 >= 40 && P2 < 50) HEX5 <= n4; 
				else if (P2 >= 50 && P2 < 60) HEX5 <= n5; 
				else if (P2 >= 60 && P2 < 70) HEX5 <= n6; 
				else if (P2 >= 70 && P2 < 80) HEX5 <= n7; 
				else if (P2 >= 80 && P2 < 90) HEX5 <= n8; 
				else HEX5 <= n9; 
		  end 
		  // HEX4 
		  begin 
				if (S2 == 0) HEX4 <= n0; 
				else if (S2 == 1) HEX4 <= n1; 
				else if (S2 == 2) HEX4 <= n2; 
				else if (S2 == 3) HEX4 <= n3; 
				else if (S2 == 4) HEX4 <= n4; 
				else if (S2 == 5) HEX4 <= n5; 
				else if (S2 == 6) HEX4 <= n6; 
				else if (S2 == 7) HEX4 <= n7; 
				else if (S2 == 8) HEX4 <= n8; 
				else HEX4 <= n9; 
		  end 
	 end 
endmodule 
	  
// ------------------------------------------------------ 
// SubModule: VGA Display 640x480 
// ------------------------------------------------------ 

module vga640x480( 
	 input wire VGA_CLK,       //pixel clock: 25MHz 
	 input wire [6:0] P1,      //Counter for P1 points 
	 input wire [6:0] P2,      //Counter for P2 points 
	 input wire [3:0] S1,      //Ones digit of P1 points 
	 input wire [3:0] S2,      //Ones digit of P2 points
	 input wire [23:0] color1, //Color of lightsaber 1
	 input wire [23:0] color2, //COlor of lightsaber 2
	 input wire reset,         //asynchronous reset 
	 output wire hsync,        //horizontal sync out 
	 output wire vsync,        //vertical sync out 
	 output reg [7:0] red,     //red vga output 
	 output reg [7:0] green,   //green vga output 
	 output reg [7:0] blue     //blue vga output 
	 ); 
		
	  // Characters in 60x30 pixels 
	  // Letter "P" 
	  reg [29:0] P[59:0]; 
			 
	  // Letter "L" 
	  reg [29:0] L[59:0];  
		
	  // Letter "A" 
	  reg [29:0] A[59:0]; 
		
	  // Letter "Y" 
	  reg [29:0] Y[59:0]; 
		
	  // Letter "E" 
	  reg [29:0] E[59:0]; 
		
	  // Letter "R" 
	  reg [29:0] R[59:0]; 
		
	  // Letter "1" 
	  reg [29:0] one[59:0]; 
		
	  // Letter "2" 
	  reg [29:0] two[59:0]; 
		
	  always @(posedge VGA_CLK) 
	  begin 
			if (reset) // Utilized to initialize 
			begin 
				// Initializing "P" 
				P[0] = 30'b000111111111111111111100000000; 
				P[1] = 30'b000111111111111111111100000000; 
				P[2] = 30'b000111111111111111111110000000; 
				P[3] = 30'b000111111000000001111110000000; 
				P[4] = 30'b000111111000000000111111000000; 
				P[5] = 30'b000111111000000000111111000000; 
				P[6] = 30'b000111111000000000011111100000; 
				P[7] = 30'b000111111000000000011111100000; 
				P[8] = 30'b000111111000000000001111110000; 
				P[9] = 30'b000111111000000000001111110000; 
				P[10] = 30'b000111111000000000000111111000; 
				P[11] = 30'b000111111000000000000111111000; 
				P[12] = 30'b000111111000000000000011111100; 
				P[13] = 30'b000111111000000000000011111100; 
				P[14] = 30'b000111111000000000000011111100; 
				P[15] = 30'b000111111000000000000011111100; 
				P[16] = 30'b000111111000000000000011111100; 
				P[17] = 30'b000111111000000000000111111000; 
				P[18] = 30'b000111111000000000000111111000; 
				P[19] = 30'b000111111000000000001111110000; 
				P[20] = 30'b000111111000000000001111110000; 
				P[21] = 30'b000111111000000000011111100000; 
				P[22] = 30'b000111111000000000011111100000; 
				P[23] = 30'b000111111000000000111111000000; 
				P[24] = 30'b000111111000000000111111000000; 
				P[25] = 30'b000111111000000001111110000000; 
				P[26] = 30'b000111111000000001111110000000; 
				P[27] = 30'b000111111111111111111110000000; 
				P[28] = 30'b000111111111111111111100000000; 
				P[29] = 30'b000111111111111111111100000000; 
				P[30] = 30'b000111111000000000000000000000; 
				P[31] = 30'b000111111000000000000000000000; 
				P[32] = 30'b000111111000000000000000000000; 
				P[33] = 30'b000111111000000000000000000000; 
				P[34] = 30'b000111111000000000000000000000; 
				P[35] = 30'b000111111000000000000000000000; 
				P[36] = 30'b000111111000000000000000000000; 
				P[37] = 30'b000111111000000000000000000000; 
				P[38] = 30'b000111111000000000000000000000; 
				P[39] = 30'b000111111000000000000000000000; 
				P[40] = 30'b000111111000000000000000000000; 
				P[41] = 30'b000111111000000000000000000000; 
				P[42] = 30'b000111111000000000000000000000; 
				P[43] = 30'b000111111000000000000000000000; 
				P[44] = 30'b000111111000000000000000000000; 
				P[45] = 30'b000111111000000000000000000000; 
				P[46] = 30'b000111111000000000000000000000; 
				P[47] = 30'b000111111000000000000000000000; 
				P[48] = 30'b000111111000000000000000000000; 
				P[49] = 30'b000111111000000000000000000000; 
				P[50] = 30'b000111111000000000000000000000; 
				P[51] = 30'b000111111000000000000000000000; 
				P[52] = 30'b000111111000000000000000000000; 
				P[53] = 30'b000111111000000000000000000000; 
				P[54] = 30'b000111111000000000000000000000; 
				P[55] = 30'b000111111000000000000000000000; 
				P[56] = 30'b000111111000000000000000000000; 
				P[57] = 30'b000111111000000000000000000000; 
				P[58] = 30'b000111111000000000000000000000; 
				P[59] = 30'b000111111000000000000000000000; 

				// Initializing "L" 
				L[0] = 30'b000111111110000000000000000000; 
				L[1] = 30'b000111111110000000000000000000; 
				L[2] = 30'b000111111110000000000000000000; 
				L[3] = 30'b000111111110000000000000000000; 
				L[4] = 30'b000111111110000000000000000000; 
				L[5] = 30'b000111111110000000000000000000; 
				L[6] = 30'b000111111110000000000000000000; 
				L[7] = 30'b000111111110000000000000000000; 
				L[8] = 30'b000111111110000000000000000000; 
				L[9] = 30'b000111111110000000000000000000; 
				L[10] = 30'b000111111110000000000000000000; 
				L[11] = 30'b000111111110000000000000000000; 
				L[12] = 30'b000111111110000000000000000000; 
				L[13] = 30'b000111111110000000000000000000; 
				L[14] = 30'b000111111110000000000000000000; 
				L[15] = 30'b000111111110000000000000000000; 
				L[16] = 30'b000111111110000000000000000000; 
				L[17] = 30'b000111111110000000000000000000; 
				L[18] = 30'b000111111110000000000000000000; 
				L[19] = 30'b000111111110000000000000000000; 
				L[20] = 30'b000111111110000000000000000000; 
				L[21] = 30'b000111111110000000000000000000; 
				L[22] = 30'b000111111110000000000000000000; 
				L[23] = 30'b000111111110000000000000000000; 
				L[24] = 30'b000111111110000000000000000000; 
				L[25] = 30'b000111111110000000000000000000; 
				L[26] = 30'b000111111110000000000000000000; 
				L[27] = 30'b000111111110000000000000000000; 
				L[28] = 30'b000111111110000000000000000000; 
				L[29] = 30'b000111111110000000000000000000; 
				L[30] = 30'b000111111110000000000000000000; 
				L[31] = 30'b000111111110000000000000000000; 
				L[32] = 30'b000111111110000000000000000000; 
				L[33] = 30'b000111111110000000000000000000; 
				L[34] = 30'b000111111110000000000000000000; 
				L[35] = 30'b000111111110000000000000000000; 
				L[36] = 30'b000111111110000000000000000000; 
				L[37] = 30'b000111111110000000000000000000; 
				L[38] = 30'b000111111110000000000000000000; 
				L[39] = 30'b000111111110000000000000000000; 
				L[40] = 30'b000111111110000000000000000000; 
				L[41] = 30'b000111111110000000000000000000; 
				L[42] = 30'b000111111110000000000000000000; 
				L[43] = 30'b000111111110000000000000000000; 
				L[44] = 30'b000111111110000000000000000000; 
				L[45] = 30'b000111111110000000000000000000; 
				L[46] = 30'b000111111110000000000000000000; 
				L[47] = 30'b000111111110000000000000000000; 
				L[48] = 30'b000111111110000000000000000000; 
				L[49] = 30'b000111111110000000000000000000; 
				L[50] = 30'b000111111111111111111111111100; 
				L[51] = 30'b000111111111111111111111111100; 
				L[52] = 30'b000111111111111111111111111100; 
				L[53] = 30'b000111111111111111111111111100; 
				L[54] = 30'b000111111111111111111111111100; 
				L[55] = 30'b000111111111111111111111111100; 
				L[56] = 30'b000111111111111111111111111100; 
				L[57] = 30'b000111111111111111111111111100; 
				L[58] = 30'b000111111111111111111111111100; 
				L[59] = 30'b000111111111111111111111111100; 
				 
				// Initializing "A" 
				A[0] = 30'b000000000001111111100000000000; 
				A[1] = 30'b000000000001111111100000000000; 
				A[2] = 30'b000000000011111111110000000000; 
				A[3] = 30'b000000000011111111110000000000; 
				A[4] = 30'b000000000111111111111000000000; 
				A[5] = 30'b000000000111111111111000000000; 
				A[6] = 30'b000000001111110011111100000000; 
				A[7] = 30'b000000001111110011111100000000; 
				A[8] = 30'b000000001111110011111100000000; 
				A[9] = 30'b000000001111110011111100000000; 
				A[10] = 30'b000000011111100001111110000000; 
				A[11] = 30'b000000011111100001111110000000; 
				A[12] = 30'b000000011111100001111110000000; 
				A[13] = 30'b000000011111100001111110000000; 
				A[14] = 30'b000000111111000000111111000000; 
				A[15] = 30'b000000111111000000111111000000; 
				A[16] = 30'b000000111111000000111111000000; 
				A[17] = 30'b000000111111000000111111000000; 
				A[18] = 30'b000001111110000000011111100000; 
				A[19] = 30'b000001111110000000011111100000; 
				A[20] = 30'b000001111110000000011111100000; 
				A[21] = 30'b000001111110000000011111100000; 
				A[22] = 30'b000011111100000000001111110000; 
				A[23] = 30'b000011111100000000001111110000; 
				A[24] = 30'b000011111100000000001111110000; 
				A[25] = 30'b000011111100000000001111110000; 
				A[26] = 30'b000111111000000000000111111000; 
				A[27] = 30'b000111111000000000000111111000; 
				A[28] = 30'b000111111000000000000111111000; 
				A[29] = 30'b000111111000000000000111111000; 
				A[30] = 30'b000111111111111111111111111000; 
				A[31] = 30'b001111111111111111111111111100; 
				A[32] = 30'b001111111111111111111111111100; 
				A[33] = 30'b001111111111111111111111111100; 
				A[34] = 30'b001111111111111111111111111100; 
				A[35] = 30'b001111111111111111111111111100; 
				A[36] = 30'b001111111000000000000111111100; 
				A[37] = 30'b001111111000000000000111111100; 
				A[38] = 30'b001111111000000000000111111100; 
				A[39] = 30'b001111111000000000000111111100; 
				A[40] = 30'b001111111000000000000111111100; 
				A[41] = 30'b001111111000000000000111111100; 
				A[42] = 30'b001111111000000000000111111100; 
				A[43] = 30'b001111111000000000000111111100; 
				A[44] = 30'b001111111000000000000111111100; 
				A[45] = 30'b001111111000000000000111111100; 
				A[46] = 30'b001111111000000000000111111100; 
				A[47] = 30'b001111111000000000000111111100; 
				A[48] = 30'b001111111000000000000111111100; 
				A[49] = 30'b001111111000000000000111111100; 
				A[50] = 30'b001111111000000000000111111100; 
				A[51] = 30'b001111111000000000000111111100; 
				A[52] = 30'b001111111000000000000111111100; 
				A[53] = 30'b001111111000000000000111111100; 
				A[54] = 30'b001111111000000000000111111100; 
				A[55] = 30'b001111111000000000000111111100; 
				A[56] = 30'b001111111000000000000111111100; 
				A[57] = 30'b001111111000000000000111111100; 
				A[58] = 30'b001111111000000000000111111100; 
				A[59] = 30'b001111111000000000000111111100; 
				 
				// Initializing "Y" 
				Y[0] = 30'b001111111100000000001111111100; 
				Y[1] = 30'b001111111100000000001111111100; 
				Y[2] = 30'b001111111100000000001111111100; 
				Y[3] = 30'b001111111100000000001111111100; 
				Y[4] = 30'b000111111110000000011111111000; 
				Y[5] = 30'b000111111110000000011111111000; 
				Y[6] = 30'b000111111110000000011111111000; 
				Y[7] = 30'b000111111110000000011111111000; 
				Y[8] = 30'b000011111111000000111111110000; 
				Y[9] = 30'b000011111111000000111111110000; 
				Y[10] = 30'b000011111111000000111111110000; 
				Y[11] = 30'b000011111111000000111111110000; 
				Y[12] = 30'b000001111111100001111111100000; 
				Y[13] = 30'b000001111111100001111111100000; 
				Y[14] = 30'b000001111111100001111111100000; 
				Y[15] = 30'b000001111111100001111111100000; 
				Y[16] = 30'b000000111111110011111111000000; 
				Y[17] = 30'b000000111111110011111111000000; 
				Y[18] = 30'b000000111111110011111111000000; 
				Y[19] = 30'b000000111111110011111111000000; 
				Y[20] = 30'b000000011111111111111110000000; 
				Y[21] = 30'b000000011111111111111110000000; 
				Y[22] = 30'b000000011111111111111110000000; 
				Y[23] = 30'b000000011111111111111110000000; 
				Y[24] = 30'b000000001111111111111100000000; 
				Y[25] = 30'b000000001111111111111100000000; 
				Y[26] = 30'b000000001111111111111100000000; 
				Y[27] = 30'b000000000111111111111000000000; 
				Y[28] = 30'b000000000111111111111000000000; 
				Y[29] = 30'b000000000111111111111000000000; 
				Y[30] = 30'b000000000011111111110000000000; 
				Y[31] = 30'b000000000011111111110000000000; 
				Y[32] = 30'b000000000011111111110000000000; 
				Y[33] = 30'b000000000011111111110000000000; 
				Y[34] = 30'b000000000011111111110000000000; 
				Y[35] = 30'b000000000011111111110000000000; 
				Y[36] = 30'b000000000011111111110000000000; 
				Y[37] = 30'b000000000011111111110000000000; 
				Y[38] = 30'b000000000011111111110000000000; 
				Y[39] = 30'b000000000011111111110000000000; 
				Y[40] = 30'b000000000011111111110000000000; 
				Y[41] = 30'b000000000011111111110000000000; 
				Y[42] = 30'b000000000011111111110000000000; 
				Y[43] = 30'b000000000011111111110000000000; 
				Y[44] = 30'b000000000011111111110000000000; 
				Y[45] = 30'b000000000011111111110000000000; 
				Y[46] = 30'b000000000011111111110000000000; 
				Y[47] = 30'b000000000011111111110000000000; 
				Y[48] = 30'b000000000011111111110000000000; 
				Y[49] = 30'b000000000011111111110000000000; 
				Y[50] = 30'b000000000011111111110000000000; 
				Y[51] = 30'b000000000011111111110000000000; 
				Y[52] = 30'b000000000011111111110000000000; 
				Y[53] = 30'b000000000011111111110000000000; 
				Y[54] = 30'b000000000011111111110000000000; 
				Y[55] = 30'b000000000011111111110000000000; 
				Y[56] = 30'b000000000011111111110000000000; 
				Y[57] = 30'b000000000011111111110000000000; 
				Y[58] = 30'b000000000011111111110000000000; 
				Y[59] = 30'b000000000011111111110000000000; 

				// Initializing "E" 
				E[0] = 30'b000111111111111111111111111000; 
				E[1] = 30'b000111111111111111111111111000; 
				E[2] = 30'b000111111111111111111111111000; 
				E[3] = 30'b000111111111111111111111111000; 
				E[4] = 30'b000111111111111111111111111000; 
				E[5] = 30'b000111111111111111111111111000; 
				E[6] = 30'b000111111111111111111111111000; 
				E[7] = 30'b000111111111111111111111111000; 
				E[8] = 30'b000111111111111111111111111000; 
				E[9] = 30'b000111111111111111111111111000; 
				E[10] = 30'b000111111111100000000000000000; 
				E[11] = 30'b000111111111100000000000000000; 
				E[12] = 30'b000111111111100000000000000000; 
				E[13] = 30'b000111111111100000000000000000; 
				E[14] = 30'b000111111111100000000000000000; 
				E[15] = 30'b000111111111100000000000000000; 
				E[16] = 30'b000111111111100000000000000000; 
				E[17] = 30'b000111111111100000000000000000; 
				E[18] = 30'b000111111111100000000000000000; 
				E[19] = 30'b000111111111100000000000000000; 
				E[20] = 30'b000111111111100000000000000000; 
				E[21] = 30'b000111111111100000000000000000; 
				E[22] = 30'b000111111111100000000000000000; 
				E[23] = 30'b000111111111100000000000000000; 
				E[24] = 30'b000111111111111111111111111000; 
				E[25] = 30'b000111111111111111111111111000; 
				E[26] = 30'b000111111111111111111111111000; 
				E[27] = 30'b000111111111111111111111111000; 
				E[28] = 30'b000111111111111111111111111000; 
				E[29] = 30'b000111111111111111111111111000; 
				E[30] = 30'b000111111111111111111111111000; 
				E[31] = 30'b000111111111111111111111111000; 
				E[32] = 30'b000111111111111111111111111000; 
				E[33] = 30'b000111111111111111111111111000; 
				E[34] = 30'b000111111111100000000000000000; 
				E[35] = 30'b000111111111100000000000000000; 
				E[36] = 30'b000111111111100000000000000000; 
				E[37] = 30'b000111111111100000000000000000; 
				E[38] = 30'b000111111111100000000000000000; 
				E[39] = 30'b000111111111100000000000000000; 
				E[40] = 30'b000111111111100000000000000000; 
				E[41] = 30'b000111111111100000000000000000; 
				E[42] = 30'b000111111111100000000000000000; 
				E[43] = 30'b000111111111100000000000000000; 
				E[44] = 30'b000111111111100000000000000000; 
				E[45] = 30'b000111111111100000000000000000; 
				E[46] = 30'b000111111111100000000000000000; 
				E[47] = 30'b000111111111100000000000000000; 
				E[48] = 30'b000111111111100000000000000000; 
				E[49] = 30'b000111111111100000000000000000; 
				E[50] = 30'b000111111111111111111111111000; 
				E[51] = 30'b000111111111111111111111111000; 
				E[52] = 30'b000111111111111111111111111000; 
				E[53] = 30'b000111111111111111111111111000; 
				E[54] = 30'b000111111111111111111111111000; 
				E[55] = 30'b000111111111111111111111111000; 
				E[56] = 30'b000111111111111111111111111000; 
				E[57] = 30'b000111111111111111111111111000; 
				E[58] = 30'b000111111111111111111111111000; 
				E[59] = 30'b000111111111111111111111111000; 
				 
				// Initializing "R" 
				R[0] = 30'b000111111111111111110000000000; 
				R[1] = 30'b000111111111111111111000000000; 
				R[2] = 30'b000111111111111111111100000000; 
				R[3] = 30'b000111111111111111111100000000; 
				R[4] = 30'b000111111111111111111110000000; 
				R[5] = 30'b000111111110000111111110000000; 
				R[6] = 30'b000111111110000011111111000000; 
				R[7] = 30'b000111111110000011111111000000; 
				R[8] = 30'b000111111110000001111111100000; 
				R[9] = 30'b000111111110000001111111100000; 
				R[10] = 30'b000111111110000000111111110000; 
				R[11] = 30'b000111111110000000111111110000; 
				R[12] = 30'b000111111110000000011111111000; 
				R[13] = 30'b000111111110000000011111111000; 
				R[14] = 30'b000111111110000000001111111100; 
				R[15] = 30'b000111111110000000001111111100; 
				R[16] = 30'b000111111110000000001111111100; 
				R[17] = 30'b000111111110000000011111111000; 
				R[18] = 30'b000111111110000000011111111000; 
				R[19] = 30'b000111111110000000111111110000; 
				R[20] = 30'b000111111110000000111111110000; 
				R[21] = 30'b000111111110000001111111100000; 
				R[22] = 30'b000111111110000001111111100000; 
				R[23] = 30'b000111111110000011111111000000; 
				R[24] = 30'b000111111110000011111111000000; 
				R[25] = 30'b000111111110000111111110000000; 
				R[26] = 30'b000111111110000111111110000000; 
				R[27] = 30'b000111111110001111111100000000; 
				R[28] = 30'b000111111111111111111100000000; 
				R[29] = 30'b000111111111111111111000000000; 
				R[30] = 30'b000111111111111111110000000000; 
				R[31] = 30'b000111111111111111100000000000; 
				R[32] = 30'b000111111111111111100000000000; 
				R[33] = 30'b000111111110111111110000000000; 
				R[34] = 30'b000111111110111111110000000000; 
				R[35] = 30'b000111111110111111110000000000; 
				R[36] = 30'b000111111110011111111000000000; 
				R[37] = 30'b000111111110011111111000000000; 
				R[38] = 30'b000111111110011111111000000000; 
				R[39] = 30'b000111111110001111111100000000; 
				R[40] = 30'b000111111110001111111100000000; 
				R[41] = 30'b000111111110001111111100000000; 
				R[42] = 30'b000111111110000111111110000000; 
				R[43] = 30'b000111111110000111111110000000; 
				R[44] = 30'b000111111110000111111110000000; 
				R[45] = 30'b000111111110000011111111000000; 
				R[46] = 30'b000111111110000011111111000000; 
				R[47] = 30'b000111111110000011111111000000; 
				R[48] = 30'b000111111110000001111111100000; 
				R[49] = 30'b000111111110000001111111100000; 
				R[50] = 30'b000111111110000001111111100000; 
				R[51] = 30'b000111111110000000111111110000; 
				R[52] = 30'b000111111110000000111111110000; 
				R[53] = 30'b000111111110000000111111110000; 
				R[54] = 30'b000111111110000000011111111000; 
				R[55] = 30'b000111111110000000011111111000; 
				R[56] = 30'b000111111110000000011111111000; 
				R[57] = 30'b000111111110000000001111111100; 
				R[58] = 30'b000111111110000000001111111100; 
				R[59] = 30'b000111111110000000001111111100; 
				 
				// Initializing "1" 
				one[0] = 30'b000000000000000001111111111000; 
				one[1] = 30'b000000000000000011111111111000; 
				one[2] = 30'b000000000000000111111111111000; 
				one[3] = 30'b000000000000001111111111111000; 
				one[4] = 30'b000000000000011111111111111000; 
				one[5] = 30'b000000000000111111111111111000; 
				one[6] = 30'b000000000001111111111111111000; 
				one[7] = 30'b000000000011111111011111111000; 
				one[8] = 30'b000000000111111110011111111000; 
				one[9] = 30'b000000001111111100011111111000; 
				one[10] = 30'b000000011111111000011111111000; 
				one[11] = 30'b000000111111110000011111111000; 
				one[12] = 30'b000000000000000000011111111000; 
				one[13] = 30'b000000000000000000011111111000; 
				one[14] = 30'b000000000000000000011111111000; 
				one[15] = 30'b000000000000000000011111111000; 
				one[16] = 30'b000000000000000000011111111000; 
				one[17] = 30'b000000000000000000011111111000; 
				one[18] = 30'b000000000000000000011111111000; 
				one[19] = 30'b000000000000000000011111111000; 
				one[20] = 30'b000000000000000000011111111000; 
				one[21] = 30'b000000000000000000011111111000; 
				one[22] = 30'b000000000000000000011111111000; 
				one[23] = 30'b000000000000000000011111111000; 
				one[24] = 30'b000000000000000000011111111000; 
				one[25] = 30'b000000000000000000011111111000; 
				one[26] = 30'b000000000000000000011111111000; 
				one[27] = 30'b000000000000000000011111111000; 
				one[28] = 30'b000000000000000000011111111000; 
				one[29] = 30'b000000000000000000011111111000; 
				one[30] = 30'b000000000000000000011111111000; 
				one[31] = 30'b000000000000000000011111111000; 
				one[32] = 30'b000000000000000000011111111000; 
				one[33] = 30'b000000000000000000011111111000; 
				one[34] = 30'b000000000000000000011111111000; 
				one[35] = 30'b000000000000000000011111111000; 
				one[36] = 30'b000000000000000000011111111000; 
				one[37] = 30'b000000000000000000011111111000; 
				one[38] = 30'b000000000000000000011111111000; 
				one[39] = 30'b000000000000000000011111111000; 
				one[40] = 30'b000000000000000000011111111000; 
				one[41] = 30'b000000000000000000011111111000; 
				one[42] = 30'b000000000000000000011111111000; 
				one[43] = 30'b000000000000000000011111111000; 
				one[44] = 30'b000000000000000000011111111000; 
				one[45] = 30'b000000000000000000011111111000; 
				one[46] = 30'b000000000000000000011111111000; 
				one[47] = 30'b000000000000000000011111111000; 
				one[48] = 30'b000000000000000000011111111000; 
				one[49] = 30'b000000000000000000011111111000; 
				one[50] = 30'b000000000000000000011111111000; 
				one[51] = 30'b000000000000000000011111111000; 
				one[52] = 30'b000000000000000000011111111000; 
				one[53] = 30'b000000000000000000011111111000; 
				one[54] = 30'b000000000000000000011111111000; 
				one[55] = 30'b000000000000000000011111111000; 
				one[56] = 30'b000000000000000000011111111000; 
				one[57] = 30'b000000000000000000011111111000; 
				one[58] = 30'b000000000000000000011111111000; 
				one[59] = 30'b000000000000000000011111111000; 

				// Initializing "2" 
				two[0] = 30'b000000011111111111110000000000; 
				two[1] = 30'b000000011111111111110000000000; 
				two[2] = 30'b000000011111111111110000000000; 
				two[3] = 30'b000000111111111111111000000000; 
				two[4] = 30'b000000111111111111111000000000; 
				two[5] = 30'b000000111111111111111000000000; 
				two[6] = 30'b000001111111111111111100000000; 
				two[7] = 30'b000001111111101111111100000000; 
				two[8] = 30'b000001111111101111111100000000; 
				two[9] = 30'b000011111111000111111110000000; 
				two[10] = 30'b000011111111000111111110000000; 
				two[11] = 30'b000011111111000111111110000000; 
				two[12] = 30'b000111111110000011111111000000; 
				two[13] = 30'b000111111110000011111111000000; 
				two[14] = 30'b000111111110000011111111000000; 
				two[15] = 30'b001111111100000001111111100000; 
				two[16] = 30'b001111111100000001111111100000; 
				two[17] = 30'b001111111100000001111111100000; 
				two[18] = 30'b001111111000000000111111110000; 
				two[19] = 30'b001111111000000000111111110000; 
				two[20] = 30'b000000000000000000011111110000; 
				two[21] = 30'b000000000000000000011111110000; 
				two[22] = 30'b000000000000000000011111110000; 
				two[23] = 30'b000000000000000000111111110000; 
				two[24] = 30'b000000000000000000111111110000; 
				two[25] = 30'b000000000000000001111111100000; 
				two[26] = 30'b000000000000000001111111100000; 
				two[27] = 30'b000000000000000011111111000000; 
				two[28] = 30'b000000000000000011111111000000; 
				two[29] = 30'b000000000000000111111110000000; 
				two[30] = 30'b000000000000000111111110000000; 
				two[31] = 30'b000000000000001111111100000000; 
				two[32] = 30'b000000000000001111111100000000; 
				two[33] = 30'b000000000000011111111000000000; 
				two[34] = 30'b000000000000011111111000000000; 
				two[35] = 30'b000000000000111111110000000000; 
				two[36] = 30'b000000000000111111110000000000; 
				two[37] = 30'b000000000001111111100000000000; 
				two[38] = 30'b000000000001111111100000000000; 
				two[39] = 30'b000000000011111111000000000000; 
				two[40] = 30'b000000000011111111000000000000; 
				two[41] = 30'b000000000111111110000000000000; 
				two[42] = 30'b000000000111111110000000000000; 
				two[43] = 30'b000000001111111100000000000000; 
				two[44] = 30'b000000001111111100000000000000; 
				two[45] = 30'b000000011111111000000000000000; 
				two[46] = 30'b000000011111111000000000000000; 
				two[47] = 30'b000000111111110000000000000000; 
				two[48] = 30'b000000111111110000000000000000; 
				two[49] = 30'b000001111111100000000000000000; 
				two[50] = 30'b000001111111100000000000000000; 
				two[51] = 30'b000011111111000000000000000000; 
				two[52] = 30'b000011111111000000000000000000; 
				two[53] = 30'b000111111110000000000000000000; 
				two[54] = 30'b000111111110000000000000000000; 
				two[55] = 30'b000111111111111111111111111000; 
				two[56] = 30'b000111111111111111111111111000; 
				two[57] = 30'b000111111111111111111111111000; 
				two[58] = 30'b000111111111111111111111111000; 
				two[59] = 30'b000111111111111111111111111000; 
			end 
	  end 
		
	 // video structure constants 
	 parameter hpixels = 800;    // horizontal pixels per line 
	 parameter vlines = 525;     // vertical lines per frame 
	 parameter hpulse = 96;    // hsync pulse length 
	 parameter vpulse = 2;     // vsync pulse length 
	 parameter hbp = 144;         // end of horizontal back porch 
	 parameter hfp = 784;         // beginning of horizontal front porch 
	 parameter vbp = 31;       // end of vertical back porch 
	 parameter vfp = 511;         // beginning of vertical front porch 
	 // active horizontal video is therefore: 784 - 144 = 640 
	 // active vertical video is therefore: 511 - 31 = 480 
		
	 // Storing the horizontal & vertical counters 
	 reg [9:0] hc; 
	 reg [9:0] vc; 

	 // Horizontal & vertical counters -- 
	 // this is how we keep track of where we are on the screen 
	 always @(posedge VGA_CLK) 
	 begin 
		  // reset condition 
		  if (reset) 
		  begin 
				hc <= 0; 
				vc <= 0; 
		  end 
		  else 
		  begin 
				// keep counting until the end of the line 
				if (hc < hpixels - 1) 
					 hc <= hc + 1; 
				else 
				// When we hit the end of the line, reset the horizontal 
				// counter and increment the vertical counter. 
				// If vertical counter is at the end of the frame, then 
				// reset that one too. 
				begin 
					 hc <= 0; 
					 if (vc < vlines - 1) 
						  vc <= vc + 1; 
					 else 
						  vc <= 0; 
				end 
				 
		  end 
	 end 
		
	 // generate sync pulses (active low) based on the  
	  // Horizontal and Vertical Counter 
	 assign hsync = (hc < hpulse) ? 0:1; 
	 assign vsync = (vc < vpulse) ? 0:1; 
		
	 always @* 
	 begin 
		  //-------------- 
		  // ROWS 0 - 60 
		  //-------------- 
		  if (vc >= vbp && vc < (vbp+60)) 
		  begin 
				if (hc >= hbp && hc < (hbp+315)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end 
				else if (hc >= (hbp+315) && hc < (hbp+325))
				begin
					 red = 0;
					 green = 0;
					 blue = 0;
				end
				else if (hc >= (hbp+325) && hc < (hbp+640))
				begin
					 red = 255;
					 green = 255;
					 blue = 255;
				end
				// Outside horizontal range, display black 
				else 
				begin 
					 red = 0; 
					 green = 0; 
					 blue = 0; 
				end 
		  end 
		  //-------------- 
		  // ROWS 60 - 120 
		  //-------------- 
		  // Displaying the letters 
		  else if (vc >= (vbp+60) && vc < (vbp+120)) 
		  begin 
				// White display 
				if (hc >= hbp && hc < (hbp+40)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end 
				// Displaying "P" for P1 
				else if (hc >= (hbp+40) && hc < (hbp+70)) 
				begin 
					 if (P[vc-vbp-60][hbp-hc+70] == 0) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 0; 
						  blue = 255; 
					 end 
				end 
				// Displaying "L" for P1 
				else if (hc >= (hbp+70) && hc < (hbp+100)) 
				begin 
					 if (L[vc-vbp-60][hbp-hc+100] == 0) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 0; 
						  blue = 255; 
					 end 
				end 
				// Displaying "A" for P1 
				else if (hc >= (hbp+100) && hc < (hbp+130)) 
				begin 
					 if (A[vc-vbp-60][hbp-hc+130] == 0) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 0; 
						  blue = 255; 
					 end 
				end 
				// Displaying "Y" for P1 
				else if (hc >= (hbp+130) && hc < (hbp+160)) 
				begin 
					 if (Y[vc-vbp-60][hbp-hc+160] == 0) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 0; 
						  blue = 255; 
					 end 
				end 
				// Displaying "E" for P1 
				else if (hc >= (hbp+160) && hc < (hbp+190)) 
				begin 
					 if (E[vc-vbp-60][hbp-hc+190] == 0) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 0; 
						  blue = 255; 
					 end 
				end 
				// Displaying "R" for P1 
				else if (hc >= (hbp+190) && hc < (hbp+220)) 
				begin 
					 if (R[vc-vbp-60][hbp-hc+220] == 0) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 0; 
						  blue = 255; 
					 end 
				end 
				// Displaying "1" for P1 
				else if (hc >= (hbp+220) && hc < (hbp+250)) 
				begin 
					 if (one[vc-vbp-60][hbp-hc+250] == 0) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 0; 
						  blue = 255; 
					 end 
				end 
				// Displaying white spaces between P1 and P2 
				else if (hc >= (hbp+250) && hc < (hbp+315)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end 
				// Put a vertical black line between
				else if (hc >= (hbp+315) && hc < (hbp+325))
				begin
					 red = 0;
					 green = 0;
					 blue = 0;
				end
				else if (hc >= (hbp+325) && hc < (hbp+360))
				begin
					 red = 255;
					 green = 255;
					 blue = 255;
				end
				// Displaying "P" for P2 
				else if (hc >= (hbp+360) && hc < (hbp+390)) 
				begin 
					 if (P[vc-vbp-60][hbp-hc+390] == 0) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 0; 
						  blue = 255; 
					 end 
				end 
				// Displaying "L" for P2 
				else if (hc >= (hbp+390) && hc < (hbp+420)) 
				begin 
					 if (L[vc-vbp-60][hbp-hc+420] == 0) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 0; 
						  blue = 255; 
					 end 
				end 
				// Displaying "A" for P2 
				else if (hc >= (hbp+420) && hc < (hbp+450)) 
				begin 
					 if (A[vc-vbp-60][hbp-hc+450] == 0) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 0; 
						  blue = 255; 
					 end 
				end 
				// Displaying "Y" for P2 
				else if (hc >= (hbp+450) && hc < (hbp+480)) 
				begin 
					 if (Y[vc-vbp-60][hbp-hc+480] == 0) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 0; 
						  blue = 255; 
					 end 
				end 
				// Displaying "E" for P2 
				else if (hc >= (hbp+480) && hc < (hbp+510)) 
				begin 
					 if (E[vc-vbp-60][hbp-hc+510] == 0) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 0; 
						  blue = 255; 
					 end 
				end 
				// Displaying "R" for P2 
				else if (hc >= (hbp+510) && hc < (hbp+540)) 
				begin 
					 if (R[vc-vbp-60][hbp-hc+540] == 0) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 0; 
						  blue = 255; 
					 end 
				end 
				// Displaying "2" for P2 
				else if (hc >= (hbp+540) && hc < (hbp+570)) 
				begin 
					 if (two[vc-vbp-60][hbp-hc+570] == 0) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 0; 
						  blue = 255; 
					 end 
				end 
				// White for the remaining pixels 
				else if (hc >= (hbp+540) && hc < (hbp+640)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end 
				// Outside horizontal range, display black 
				else 
				begin 
					 red = 0; 
					 green = 0; 
					 blue = 0; 
				end 
		  end 
		  //--------------- 
		  // ROWS 120 - 170 
		  //--------------- 
		  // Display more white to make difference
		  else if (vc >= (vbp+120) && vc < (vbp+170)) 
		  begin 
				// Display all white 
				if (hc >= hbp && hc < (hbp+315)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end 
				// Put a vertical black line between
				else if (hc >= (hbp+315) && hc < (hbp+325))
				begin
					 red = 0;
					 green = 0;
					 blue = 0;
				end
				else if (hc >= (hbp+325) && hc < (hbp+640))
				begin
					 red = 255;
					 green = 255;
					 blue = 255;
				end
				// Outside horizontal range, display black 
				else 
				begin 
					 red = 0; 
					 green = 0; 
					 blue = 0; 
				end 
		  end 
		  //--------------- 
		  // ROWS 170 - 175 
		  //--------------- 
		  // Display the top part of 2nd hilt
		  else if (vc >= (vbp+170) && vc < (vbp+175)) 
		  begin 
				// Display White 
				if (hc >= hbp && hc < (hbp+315)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end
				// Black line separator
				else if (hc >= (hbp+315) && hc < (hbp+325))
				begin
					 red = 0;
					 green = 0;
					 blue = 0;
				end
				else if (hc >= (hbp+325) && hc < (hbp+600))
				begin
					 red = 255;
					 green = 255;
					 blue = 255;
				end
				// Put Black part of the hilt
				else if (hc >= (hbp+600) && hc < (hbp+610))
				begin
					 red = 0;
					 green = 0;
					 blue = 0;
				end
				else if (hc >= (hbp+610) && hc < (hbp+640))
				begin
					 red = 255;
					 green = 255;
					 blue = 255;
				end
				// Outside horizontal range, display black 
				else 
				begin 
					 red = 0; 
					 green = 0; 
					 blue = 0; 
				end 
		  end 
		  //--------------- 
		  // ROWS 175 - 180 
		  //---------------
		  else if (vc >= (vbp+175) && vc < (vbp+180))
		  begin
				// Lower part of Hilt 1
				if (hc >= hbp && hc < (hbp+20))
				begin
					red = 192;
					green = 192;
					blue = 192;
				end
				// Display white for the rest
				else if (hc >= (hbp+20) && hc < (hbp+315))
				begin
					red = 255;
					green = 255;
					blue = 255;
				end
				// Black line split
				else if (hc >= (hbp+315) && hc < (hbp+325))
				begin
					red = 0;
					green = 0;
					blue = 0;
				end
				else if (hc >= (hbp+325) && hc < (hbp+570))
				begin
					red = 255;
					green = 255;
					blue = 255;
				end
				else if (hc >= (hbp+570) && hc < (hbp+580))
				begin
					red = 0;
					green = 0;
					blue = 0;
				end
				else if (hc >= (hbp+580) && hc < (hbp+600))
				begin
					red = 255;
					green = 255;
					blue = 255;
				end
				else if (hc >= (hbp+600) && hc < (hbp+610))
				begin
					red = 0;
					green = 0;
					blue = 0;
				end
				else if (hc >= (hbp+610) && hc < (hbp+615))
				begin
					red = 255;
					green = 255;
					blue = 255;
				end
				else if (hc >= (hbp+615) && hc < (hbp+640))
				begin
					red = 0;
					green = 0;
					blue = 0;
				end
				// Gone out of range
				else
				begin
					red = 0;
					green = 0;
					blue = 0;
				end
		  end
		  //--------------- 
		  // ROWS 180 - 210 
		  //---------------
		  // Bulk of the hilt and color of the blade
		  else if (vc >= (vbp+180) && vc < (vbp+210))
		  begin
				if (hc >= hbp && hc < (hbp+25))
				begin
					red = 192;
					green = 192;
					blue = 192;
				end
				else if (hc >= (hbp+25) && hc < (hbp+70))
				begin
					red = 224;
					green = 224;
					blue = 224;
				end
				// Lightsaber COlor 1
				else if (hc >= (hbp+70) && hc < (hbp+315))
				begin
					red = color1[23:16];
					green = color1[15:8];
					blue = color1[7:0];
				end
				// Black line separator
				else if (hc >= (hbp+315) && hc < (hbp+325))
				begin
					red = 0;
					green = 0;
					blue = 0;
				end
				// Lightsaber Color 2
				else if (hc >= (hbp+325) && hc < (hbp+570))
				begin
					red = color2[23:16];
					green = color2[15:8];
					blue = color2[7:0];
				end
				else if (hc >= (hbp+570) && hc < (hbp+580))
				begin
					red = 0;
					green = 0;
					blue = 0;
				end
				else if (hc >= (hbp+580) && hc < (hbp+600))
				begin
					red = 32;
					green = 32;
					blue = 32;
				end
				else if (hc >= (hbp+600) && hc < (hbp+610))
				begin
					red = 0;
					green = 0;
					blue = 0;
				end
				else if (hc >= (hbp+610) && hc < (hbp+615))
				begin
					red = 32;
					green = 32;
					blue = 32;
				end
				else if (hc >= (hbp+615) && hc < (hbp+640))
				begin
					red = 0;
					green = 0;
					blue = 0;
				end
				// At the end of vertical range
				else
				begin
					red = 0;
					green = 0;
					blue = 0;
				end
		  end
		  //--------------- 
		  // ROWS 210 - 215 
		  //---------------
		  else if (vc >= (vbp+210) && vc < (vbp+215))
		  begin
				// Part of Hilt 1
				if (hc >= hbp && hc < (hbp+20))
				begin
					red = 192;
					green = 192;
					blue = 192;
				end
				else if (hc >= (hbp+20) && hc < (hbp+52))
				begin
					red = 255;
					green = 255;
					blue = 255;
				end
				else if (hc >= (hbp+52) && hc < (hbp+57))
				begin
					red = 205;
					green = 205;
					blue = 205;
				end
				else if (hc >= (hbp+57) && hc < (hbp+62))
				begin
					red = 255;
					green = 255;
					blue = 255;
				end
				else if (hc >= (hbp+62) && hc < (hbp+67))
				begin
					red = 205;
					green = 205;
					blue = 205;
				end
				else if (hc >= (hbp+67) && hc < (hbp+315))
				begin
					red = 255;
					green = 255;
					blue = 255;
				end
				// Black line split
				else if (hc >= (hbp+315) && hc < (hbp+325))
				begin
					red = 0;
					green = 0;
					blue = 0;
				end
				else if (hc >= (hbp+325) && hc < (hbp+570))
				begin
					red = 255;
					green = 255;
					blue = 255;
				end
				else if (hc >= (hbp+570) && hc < (hbp+580))
				begin
					red = 0;
					green = 0;
					blue = 0;
				end
				else if (hc >= (hbp+580) && hc < (hbp+615))
				begin
					red = 255;
					green = 255;
					blue = 255;
				end
				else if (hc >= (hbp+615) && hc < (hbp+640))
				begin
					red = 0;
					green = 0;
					blue = 0;
				end
				// Reached end of vertical range
				else
				begin
					red = 0;
					green = 0;
					blue = 0;
				end
		  end
		  //--------------- 
		  // ROWS 215 - 220 
		  //---------------
		  else if (vc >= (vbp+215) && vc < (vbp+220))
		  begin
				if (hc >= hbp && hc < (hbp+62))
				begin
					red = 255;
					green = 255;
					blue = 255;
				end
				else if (hc >= (hbp+62) && hc < (hbp+67))
				begin
					red = 205;
					green = 205;
					blue = 205;
				end
				else if (hc >= (hbp+67) && hc < (hbp+315))
				begin
					red = 255;
					green = 255;
					blue = 255;
				end
				// Put a vertical black line between
				else if (hc >= (hbp+315) && hc < (hbp+325))
				begin
					 red = 0;
					 green = 0;
					 blue = 0;
				end
				else if (hc >= (hbp+325) && hc < (hbp+640))
				begin
					 red = 255;
					 green = 255;
					 blue = 255;
				end
				// Reached end of range
				else
				begin
					red = 0;
					green = 0;
					blue = 0;
				end
		  end
		  //--------------- 
		  // ROWS 220 - 240 
		  //--------------- 
		  // Display more white 
		  else if (vc >= (vbp+220) && vc < (vbp+240)) 
		  begin 
				if (hc >= hbp && hc < (hbp+315)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end 
				// Put a vertical black line between
				else if (hc >= (hbp+315) && hc < (hbp+325))
				begin
					 red = 0;
					 green = 0;
					 blue = 0;
				end
				else if (hc >= (hbp+325) && hc < (hbp+640))
				begin
					 red = 255;
					 green = 255;
					 blue = 255;
				end
				else 
				begin 
					 red = 0; 
					 green = 0; 
					 blue = 0; 
				end 
		  end 
			
		  //------------------------------------------------------------- 
		  // NUMBERS DISPLAY STARTS BELOW (Will be difficult) 
		  //------------------------------------------------------------- 
			
		  //--------------- 
		  // ROWS 240 - 265 
		  //--------------- 
		  else if (vc >= (vbp+240) && vc < (vbp+265)) 
		  begin 
				// White in the first few. 
				if (hc >= hbp && hc < (hbp+40)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end 
				// -------------------------------- 
				// Tens digit of Player 1 
				// -------------------------------- 
				// ---------------- 
				// Zone 1 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+40) && hc < (hbp+65)) 
				begin 
					 if (P1 >= 10 && P1 < 20) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// ---------------- 
				// Zone 2 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+65) && hc < (hbp+115)) 
				begin 
					 if ((P1 >= 10 && P1 < 20) | 
						  (P1 >= 40 && P1 < 50)) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// ---------------- 
				// Zone 3 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+115) && hc < (hbp+140)) 
				begin 
					 red = 0; 
					 green = 153; 
					 blue = 0; 
				end 
				// Whiteness to make space 
				else if (hc >= (hbp+140) && hc < (hbp+180)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end 
				// -------------------------------- 
				// Ones digit of Player 1 
				// -------------------------------- 
				else if (hc >= (hbp+180) && hc < (hbp+205)) 
				begin 
				// ---------------- 
				// Zone 1 of number (Copy and Paste) 
				// ---------------- 
					 if (S1 == 1) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// ---------------- 
				// Zone 2 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+205) && hc < (hbp+255)) 
				begin 
					 if ((S1 == 1) | 
						  (S1 == 4)) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// ---------------- 
				// Zone 3 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+255) && hc < (hbp+280)) 
				begin 
					 red = 0; 
					 green = 153; 
					 blue = 0; 
				end 
				// Whiteness to make space 
				else if (hc >= (hbp+280) && hc < (hbp+315)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end 
				// Put a vertical black line between
				else if (hc >= (hbp+315) && hc < (hbp+325))
				begin
					 red = 0;
					 green = 0;
					 blue = 0;
				end
				else if (hc >= (hbp+325) && hc < (hbp+360))
				begin
					 red = 255;
					 green = 255;
					 blue = 255;
				end
				// -------------------------------- 
				// Tens digit of Player 2 
				// -------------------------------- 
				// ---------------- 
				// Zone 1 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+360) && hc < (hbp+385)) 
				begin 
					 if (P2 >= 10 && P2 < 20) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// ---------------- 
				// Zone 2 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+385) && hc < (hbp+435)) 
				begin 
					 if ((P2 >= 10 && P2 < 20) | 
						  (P2 >= 40 && P2 < 50)) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// ---------------- 
				// Zone 3 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+435) && hc < (hbp+460)) 
				begin 
					 red = 0; 
					 green = 153; 
					 blue = 0; 
				end 
				// Whiteness to make space 
				else if (hc >= (hbp+460) && hc < (hbp+500)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end 
				// -------------------------------- 
				// Ones digit of Player 2 
				// -------------------------------- 
				// ---------------- 
				// Zone 1 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+500) && hc < (hbp+525)) 
				begin 
					 if (S2 == 1) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// ---------------- 
				// Zone 2 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+525) && hc < (hbp+575)) 
				begin 
					 if ((S2 == 1) | 
						  (S2 == 4)) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// ---------------- 
				// Zone 3 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+575) && hc < (hbp+600)) 
				begin 
					 red = 0; 
					 green = 153; 
					 blue = 0; 
				end 
				// Whiteness to make space 
				else if (hc >= (hbp+600) && hc < (hbp+640)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end 
				// Gone out of range now. 
				else 
				begin 
					 red = 0; 
					 green = 0; 
					 blue = 0; 
				end 
		  end 
		  //--------------- 
		  // ROWS 265 - 325 
		  //--------------- 
		  else if (vc >= (vbp+265) && vc < (vbp+325)) 
		  begin 
				// White in the first few. 
				if (hc >= hbp && hc < (hbp+40)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end 
				// -------------------------------- 
				// Tens digit of Player 1 
				// -------------------------------- 
				// ---------------- 
				// Zone 1 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+40) && hc < (hbp+65)) 
				begin 
					 if ((P1 >= 10 && P1 < 40) | 
						  (P1 >= 70 && P1 < 80)) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// ---------------- 
				// Zone 2 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+65) && hc < (hbp+115)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end 
				// ---------------- 
				// Zone 3 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+115) && hc < (hbp+140)) 
				begin 
					 if (P1 >= 50 && P1 < 70) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// Whiteness to make space 
				else if (hc >= (hbp+140) && hc < (hbp+180)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end 
				// -------------------------------- 
				// Ones digit of Player 1 
				// -------------------------------- 
				// ---------------- 
				// Zone 1 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+180) && hc < (hbp+205)) 
				begin 
					 if ((S1 >= 1 && S1 < 4) | 
						  (S1 == 7)) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// ---------------- 
				// Zone 2 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+205) && hc < (hbp+255)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end 
				// ---------------- 
				// Zone 3 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+255) && hc < (hbp+280)) 
				begin 
				if (S1 >= 5 && S1 < 7) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// Whiteness to make space 
				else if (hc >= (hbp+280) && hc < (hbp+315)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end 
				// Put a vertical black line between
				else if (hc >= (hbp+315) && hc < (hbp+325))
				begin
					 red = 0;
					 green = 0;
					 blue = 0;
				end
				else if (hc >= (hbp+325) && hc < (hbp+360))
				begin
					 red = 255;
					 green = 255;
					 blue = 255;
				end 
				// -------------------------------- 
				// Tens digit of Player 2 
				// -------------------------------- 
				// ---------------- 
				// Zone 1 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+360) && hc < (hbp+385)) 
				begin 
					 if ((P2 >= 10 && P2 < 40) | 
						  (P2 >= 70 && P2 < 80)) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// ---------------- 
				// Zone 2 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+385) && hc < (hbp+435)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end 
				// ---------------- 
				// Zone 3 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+435) && hc < (hbp+460)) 
				begin 
				if (P2 >= 50 && P2 < 70) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// Whiteness to make space 
				else if (hc >= (hbp+460) && hc < (hbp+500)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end 
				// -------------------------------- 
				// Ones digit of Player 2 
				// -------------------------------- 
				// ---------------- 
				// Zone 1 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+500) && hc < (hbp+525)) 
				begin 
					 if ((S2 >= 1 && S2 < 4) | 
						  (S2 == 7)) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// ---------------- 
				// Zone 2 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+525) && hc < (hbp+575)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end 
				// ---------------- 
				// Zone 3 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+575) && hc < (hbp+600)) 
				begin 
				if (S2 >= 5 && S2 < 7) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// Whiteness to make space 
				else if (hc >= (hbp+600) && hc < (hbp+640)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end 
				// Gone out of range now. 
				else 
				begin 
					 red = 0; 
					 green = 0; 
					 blue = 0; 
				end 
		  end 
		  //--------------- 
		  // ROWS 325 - 355 
		  //--------------- 
		  else if (vc >= (vbp+325) && vc < (vbp+355)) 
		  begin 
				// White in the first few. 
				if (hc >= hbp && hc < (hbp+40)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end 
				// -------------------------------- 
				// Tens digit of Player 1 
				// -------------------------------- 
				// ---------------- 
				// Zone 1 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+40) && hc < (hbp+65)) 
				begin 
					 if ((P1 >= 10 && P1 < 20) | 
						  (P1 >= 70 && P1 < 80)) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// ---------------- 
				// Zone 2 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+65) && hc < (hbp+115)) 
				begin 
					 if ((P1 >= 0 && P1 < 20) | 
						  (P1 >= 70 && P1 < 80)) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// ---------------- 
				// Zone 3 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+115) && hc < (hbp+140)) 
				begin 
					 red = 0; 
					 green = 153; 
					 blue = 0; 
				end 
				// Whiteness to make space 
				else if (hc >= (hbp+140) && hc < (hbp+180)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end 
				// -------------------------------- 
				// Ones digit of Player 1 
				// -------------------------------- 
				// ---------------- 
				// Zone 1 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+180) && hc < (hbp+205)) 
				begin 
					 if ((S1 == 1) | 
						  (S1 == 7)) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// ---------------- 
				// Zone 2 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+205) && hc < (hbp+255)) 
				begin 
					 if ((S1 >= 0 && S1 < 2) | 
						  (S1 == 7)) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// ---------------- 
				// Zone 3 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+255) && hc < (hbp+280)) 
				begin 
					 red = 0; 
					 green = 153; 
					 blue = 0; 
				end 
				// Whiteness to make space 
				else if (hc >= (hbp+280) && hc < (hbp+315)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end 
				// Put a vertical black line between
				else if (hc >= (hbp+315) && hc < (hbp+325))
				begin
					 red = 0;
					 green = 0;
					 blue = 0;
				end
				else if (hc >= (hbp+325) && hc < (hbp+360))
				begin
					 red = 255;
					 green = 255;
					 blue = 255;
				end
				// -------------------------------- 
				// Tens digit of Player 2 
				// -------------------------------- 
				// ---------------- 
				// Zone 1 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+360) && hc < (hbp+385)) 
				begin 
					 if ((P2 >= 10 && P2 < 20) | 
						  (P2 >= 70 && P2 < 80)) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// ---------------- 
				// Zone 2 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+385) && hc < (hbp+435)) 
				begin 
					 if ((P2 >= 0 && P2 < 20) | 
						  (P2 >= 70 && P2 < 80)) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// ---------------- 
				// Zone 3 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+435) && hc < (hbp+460)) 
				begin 
					 red = 0; 
					 green = 153; 
					 blue = 0; 
				end 
				// Whiteness to make space 
				else if (hc >= (hbp+460) && hc < (hbp+500)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end 
				// -------------------------------- 
				// Ones digit of Player 2 
				// -------------------------------- 
				// ---------------- 
				// Zone 1 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+500) && hc < (hbp+525)) 
				begin 
					 if ((S2 == 1) | 
						  (S2 == 7)) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// ---------------- 
				// Zone 2 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+525) && hc < (hbp+575)) 
				begin 
					 if ((S2 >= 0 && S2 < 2) | 
						  (S2 == 7)) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// ---------------- 
				// Zone 3 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+575) && hc < (hbp+600)) 
				begin 
					 red = 0; 
					 green = 153; 
					 blue = 0; 
				end 
				// Whiteness to make space 
				else if (hc >= (hbp+600) && hc < (hbp+640)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end 
				// Gone out of range now. 
				else 
				begin 
					 red = 0; 
					 green = 0; 
					 blue = 0; 
				end 
		  end 
		  //--------------- 
		  // ROWS 355 - 415 
		  //--------------- 
		  else if (vc >= (vbp+355) && vc < (vbp+415)) 
		  begin 
				// White in the first few. 
				if (hc >= hbp && hc < (hbp+40)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end 
				// -------------------------------- 
				// Tens digit of Player 1 
				// -------------------------------- 
				// ---------------- 
				// Zone 1 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+40) && hc < (hbp+65)) 
				begin 
					 if ((P1 >= 10 && P1 < 20) | 
						  (P1 >= 30 && P1 < 60) | 
						  (P1 >= 70 && P1 < 80) | 
						  (P1 >= 90 && P1 < 100)) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// ---------------- 
				// Zone 2 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+65) && hc < (hbp+115)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end 
				// ---------------- 
				// Zone 3 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+115) && hc < (hbp+140)) 
				begin 
					 if (P1 >= 20 && P1 < 30) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// Whiteness to make space 
				else if (hc >= (hbp+140) && hc < (hbp+180)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end 
				// -------------------------------- 
				// Ones digit of Player 1 
				// -------------------------------- 
				// ---------------- 
				// Zone 1 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+180) && hc < (hbp+205)) 
				begin 
					 if ((S1 == 1) | 
						  (S1 >= 3 && S1 < 6) | 
						  (S1 == 7) | 
						  (S1 == 9)) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// ---------------- 
				// Zone 2 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+205) && hc < (hbp+255)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end 
				// ---------------- 
				// Zone 3 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+255) && hc < (hbp+280)) 
				begin 
					 if (S1 == 2) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// Whiteness to make space 
				else if (hc >= (hbp+280) && hc < (hbp+315)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end 
				// Put a vertical black line between
				else if (hc >= (hbp+315) && hc < (hbp+325))
				begin
					 red = 0;
					 green = 0;
					 blue = 0;
				end
				else if (hc >= (hbp+325) && hc < (hbp+360))
				begin
					 red = 255;
					 green = 255;
					 blue = 255;
				end 
				// -------------------------------- 
				// Tens digit of Player 2 
				// -------------------------------- 
				// ---------------- 
				// Zone 1 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+360) && hc < (hbp+385)) 
				begin 
					 if ((P2 >= 10 && P2 < 20) | 
						  (P2 >= 30 && P2 < 60) | 
						  (P2 >= 70 && P2 < 80) | 
						  (P2 >= 90 && P2 < 100)) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// ---------------- 
				// Zone 2 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+385) && hc < (hbp+435)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end 
				// ---------------- 
				// Zone 3 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+435) && hc < (hbp+460)) 
				begin 
					 if (P2 >= 20 && P2 < 30) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// Whiteness to make space 
				else if (hc >= (hbp+460) && hc < (hbp+500)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end 
				// -------------------------------- 
				// Ones digit of Player 2 
				// -------------------------------- 
				// ---------------- 
				// Zone 1 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+500) && hc < (hbp+525)) 
				begin 
					 if ((S2 == 1) | 
						  (S2 >= 3 && S2 < 6) | 
						  (S2 == 7) | 
						  (S2 == 9)) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// ---------------- 
				// Zone 2 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+525) && hc < (hbp+575)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end 
				// ---------------- 
				// Zone 3 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+575) && hc < (hbp+600)) 
				begin 
					 if (S2 == 2) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// Whiteness to make space 
				else if (hc >= (hbp+600) && hc < (hbp+640)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end 
				// Gone out of range now. 
				else 
				begin 
					 red = 0; 
					 green = 0; 
					 blue = 0; 
				end 
		  end 
		  //--------------- 
		  // ROWS 415 - 440 
		  //--------------- 
		  else if (vc >= (vbp+415) && vc < (vbp+440)) 
		  begin 
				// White in the first few. 
				if (hc >= hbp && hc < (hbp+40)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end 
				// -------------------------------- 
				// Tens digit of Player 1 
				// -------------------------------- 
				// ---------------- 
				// Zone 1 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+40) && hc < (hbp+65)) 
				begin 
					 if ((P1 >= 10 && P1 < 20) | 
						  (P1 >= 40 && P1 < 50) | 
						  (P1 >= 70 && P1 < 80) | 
						  (P1 >= 90 && P1 < 100)) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// ---------------- 
				// Zone 2 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+65) && hc < (hbp+115)) 
				begin 
					 if ((P1 >= 10 && P1 < 20) | 
						  (P1 >= 40 && P1 < 50) | 
						  (P1 >= 70 && P1 < 80) | 
						  (P1 >= 90 && P1 < 100)) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// ---------------- 
				// Zone 3 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+115) && hc < (hbp+140)) 
				begin 
					 red = 0; 
					 green = 153; 
					 blue = 0; 
				end 
				// Whiteness to make space 
				else if (hc >= (hbp+140) && hc < (hbp+180)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end 
				// -------------------------------- 
				// Ones digit of Player 1 
				// -------------------------------- 
				// ---------------- 
				// Zone 1 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+180) && hc < (hbp+205)) 
				begin 
					 if ((S1 == 1) | 
						  (S1 == 4) | 
						  (S1 == 7) | 
						  (S1 == 9)) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// ---------------- 
				// Zone 2 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+205) && hc < (hbp+255)) 
				begin 
					 if ((S1 == 1) | 
						  (S1 == 4) | 
						  (S1 == 7) | 
						  (S1 == 9)) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// ---------------- 
				// Zone 3 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+255) && hc < (hbp+280)) 
				begin 
					 red = 0; 
					 green = 153; 
					 blue = 0; 
				end 
				// Whiteness to make space 
				else if (hc >= (hbp+280) && hc < (hbp+315)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end 
				// Put a vertical black line between
				else if (hc >= (hbp+315) && hc < (hbp+325))
				begin
					 red = 0;
					 green = 0;
					 blue = 0;
				end
				else if (hc >= (hbp+325) && hc < (hbp+360))
				begin
					 red = 255;
					 green = 255;
					 blue = 255;
				end 
				// -------------------------------- 
				// Tens digit of Player 2 
				// -------------------------------- 
				// ---------------- 
				// Zone 1 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+360) && hc < (hbp+385)) 
				begin 
					 if ((P2 >= 10 && P2 < 20) | 
						  (P2 >= 40 && P2 < 50) | 
						  (P2 >= 70 && P2 < 80) | 
						  (P2 >= 90 && P2 < 100)) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// ---------------- 
				// Zone 2 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+385) && hc < (hbp+435)) 
				begin 
					 if ((P2 >= 10 && P2 < 20) | 
						  (P2 >= 40 && P2 < 50) | 
						  (P2 >= 70 && P2 < 80) | 
						  (P2 >= 90 && P2 < 100)) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// ---------------- 
				// Zone 3 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+435) && hc < (hbp+460)) 
				begin 
					 red = 0; 
					 green = 153; 
					 blue = 0; 
				end 
				// Whiteness to make space 
				else if (hc >= (hbp+460) && hc < (hbp+500)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end 
				// -------------------------------- 
				// Ones digit of Player 2 
				// -------------------------------- 
				// ---------------- 
				// Zone 1 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+500) && hc < (hbp+525)) 
				begin 
					 if ((S2 == 1) | 
						  (S2 == 4) | 
						  (S2 == 7) | 
						  (S2 == 9)) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// ---------------- 
				// Zone 2 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+525) && hc < (hbp+575)) 
				begin 
					 if ((S2 == 1) | 
						  (S2 == 4) | 
						  (S2 == 7) | 
						  (S2 == 9)) 
					 begin 
						  red = 255; 
						  green = 255; 
						  blue = 255; 
					 end 
					 else 
					 begin 
						  red = 0; 
						  green = 153; 
						  blue = 0; 
					 end 
				end 
				// ---------------- 
				// Zone 3 of number (Copy and Paste) 
				// ---------------- 
				else if (hc >= (hbp+575) && hc < (hbp+600)) 
				begin 
					 red = 0; 
					 green = 153; 
					 blue = 0; 
				end 
				// Whiteness to make space 
				else if (hc >= (hbp+600) && hc < (hbp+640)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end 
				// Gone out of range now. 
				else 
				begin 
					 red = 0; 
					 green = 0; 
					 blue = 0; 
				end 
		  end 
			
		  //------------------------------------------------------------- 
		  // NUMBERS DISPLAY FINISHED ABOVE 
		  //------------------------------------------------------------- 
			
		  //--------------- 
		  // ROWS 440 - 480 
		  //--------------- 
		  // Display more white 
		  else if (vc >= (vbp+440) && vc < (vbp+480)) 
		  begin 
				if (hc >= hbp && hc < (hbp+315)) 
				begin 
					 red = 255; 
					 green = 255; 
					 blue = 255; 
				end
				// Put a vertical black line between
				else if (hc >= (hbp+315) && hc < (hbp+325))
				begin
					 red = 0;
					 green = 0;
					 blue = 0;
				end
				else if (hc >= (hbp+325) && hc < (hbp+640))
				begin
					 red = 255;
					 green = 255;
					 blue = 255;
				end
				else 
				begin 
					 red = 0; 
					 green = 0; 
					 blue = 0; 
				end 
		  end 
		  //--------------- 
		  // ROWS 480+ (Outside) 
		  //--------------- 
		// we're outside active vertical range so display black 
		else 
		begin 
				red = 0; 
				green = 0; 
				blue = 0; 
		end 
	end 

endmodule 

// ------------------------------------------------------ 
// Submodule: Debouncer (Taken from EECS270 lab) 
// ------------------------------------------------------ 

module debouncer( 
	 input clk,             //this is a 50MHz clock provided on FPGA pin PIN_Y2 
	 input PB,              //this is the input to be debounced 
	 output reg PB_state //this is the debounced switch 
); 

	 // Synchronize the switch input to the clock 
	 reg PB_sync_0; 
	 always @(posedge clk) PB_sync_0 <= PB; 
	 reg PB_sync_1; 
	 always @(posedge clk) PB_sync_1 <= PB_sync_0; 

	 // Debounce the switch 
	 reg [15:0] PB_cnt; 
	 always @(posedge clk) 
		  if(PB_state==PB_sync_1) 
				 PB_cnt <= 0; 
		  else 
	 begin 
			PB_cnt <= PB_cnt + 1'b1;  
			if(PB_cnt == 16'hffff) PB_state <= ~PB_state;  
	 end 
	  
endmodule